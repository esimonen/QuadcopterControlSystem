��m o d u l e   i n e r t _ i n t f _ t b ( ) ;  
 	  
 	 l o g i c   c l k ;  
 	 l o g i c   M I S O ; 	 	 	 	 	 / /   S P I   i n p u t   f r o m   i n e r t i a l   s e n s o r  
 	 l o g i c   I N T ; 	 	 	 	 	 / /   g o e s   h i g h   w h e n   m e a s u r e m e n t   r e a d y  
 	 l o g i c   s t r t _ c a l ; 	 	 	 	 / /   f r o m   c o m a n d   c o n f i g .     I n d i c a t e s   w e   s h o u l d   s t a r t   c a l i b r a t i o n  
 	      
 	 l o g i c   [ 7 : 0 ]   L E D ;                         / /   o u t p u t   t o   L E D   a r r a y   o n   f p g a   b o a r d  
 	 l o g i c   S S _ n , S C L K , M O S I ; 	 	 / /   S P I   o u t p u t s  
  
         l o g i c   R S T _ n ;         / /   s i m u l a t e d   ' r e s e t   b u t t o n '   o n   f p g a  
         l o g i c   N E X T ;           / /   s i m u l a t e d   ' n e x t   b u t t o n '   o n   f p g a  
  
 	 S P I _ i N E M O 2   i N e m o ( . S S _ n ( S S _ n ) , . S C L K ( S C L K ) , . M I S O ( M I S O ) , . M O S I ( M O S I ) , . I N T ( I N T ) ) ;  
 	 i n e r t _ i n t f _ t e s t   i D U T ( . c l k ( c l k ) ,   . N E X T ( N E X T ) ,   . R S T _ n ( R S T _ n ) ,   . L E D ( L E D ) ,   . S S _ n ( S S _ n ) ,   . S C L K ( S C L K ) ,   . M O S I ( M O S I ) ,   . M I S O ( M I S O ) ,   . I N T ( I N T ) ) ;  
  
 	 i n i t i a l   b e g i n  
 	 	 c l k   =   0 ;  
 	 	 R S T _ n   =   1 ;  
                 N E X T   =   1 ;  
  
                 @ ( p o s e d g e   i N E M O 2 . P O R _ n ) ;   / /   w a i t   f o r   n e m o   t o   p o w e r   u p   a n d   s e t u p  
 	 	 r e p e a t   ( 2 )   @ ( p o s e d g e   c l k ) ;   R S T _ n   =   0 ;   / /   w a i t   o n   p u s h   b u t t o n ' s   r e s e t   t o   s y n c  
 	 	 r e p e a t   ( 2 )   @ ( p o s e d g e   c l k )   N E X T   =   0 ;   / /   d e a s s e r t   r e s e t  
 	 	  
 	 	 / /   c h e c k   t h a t   N E M O _ s e t u p   g e t s   a s s e r t e d   i n   a   r e a s o n a b l e   t i m e  
 	 	 f o r k  
 	 	 	 b e g i n   :   t i m e o u t  
 	 	 	 	 r e p e a t ( 2 1 0 0 0 0 ) @ ( p o s e d g e   c l k ) ;  
 	 	 	 	 $ d i s p l a y ( " E R R O R :   t i m e o u t   o u t   w a i t i n g   f o r   N E M O _ s e t u p   t o   a s s e r t " ) ;  
 	 	 	 	 $ s t o p ;  
 	 	 	 e n d  
 	 	 	 b e g i n  
 	 	 	 	 @ ( p o s e d g e   i N e m o . N E M O _ s e t u p ) ;  
 	 	 	 	 d i s a b l e   t i m e o u t ;  
 	 	 	 e n d  
 	 	 j o i n  
 	 	  
 	 	 $ s t o p ;  
 	 	  
 	 e n d  
 	  
 	 / /   c l o c k  
 	 a l w a y s  
 	 	 # 5   c l k   =   ~ c l k ;  
 e n d m o d u l e  
 